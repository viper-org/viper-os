func @PutPixel(x: i32, y: i32, color: i32) -> void;